//=========================================================================
// 5-Stage Bypass Pipelined Processor Control
//=========================================================================

`ifndef LAB2_PROC_PIPELINED_PROC_ALT_CTRL_V
`define LAB2_PROC_PIPELINED_PROC_ALT_CTRL_V

module lab2_proc_PipelinedProcAltCtrl
(
  input  logic        clk,
 input  logic        reset
);

// copy in the baseline design and start working on the alternative!

endmodule

`endif

